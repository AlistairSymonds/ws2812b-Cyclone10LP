entity ws2812Controller is



end entity;

architecture